module axi_dut (
    
);



endmodule