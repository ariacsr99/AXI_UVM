// Common macro definitions for AXI UVM testbench

// Default Clock and Reset
`define AXI_CLOCK vif.axi_tb_ACLK
`define AXI_RESET vif.axi_tb_ARESETn